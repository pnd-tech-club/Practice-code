Your current HP is:  - 6.0 
- 6.0 
rength: 6.0
Dexterity: 6.0
Constitution: 6.0
Intelligence: 6.0
Wisdom: 6.0
Charisma: 6.0
Abilities: h
Gold: 6.0
Gear: h
Max HP: 6.0
Current HP: 6.0
Level: 6.0
